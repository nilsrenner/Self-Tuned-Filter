.title Experiment 5 - VCF

* LIBRARIES
.inc tl082.cir
.inc mpy634.cir

* PARAMETER
.param Vsup=15

R1 N010 N002 1k
R2 N011 N006 2k
R3 N013 N007 1k
R4 N002 N013 1k
R5 N013 N016 1k
R6 N016 N015 1k
R7 N015 N006 64k
R8 N015 N008 500
R9 N001 N014 100k
R10 N001 N009 10
R11 N012 N005 1k

C1 N003 N010 200n
C2 N004 N011 1u
C3 N009 N012 100n

* OPAMPs
XU1 0 N010 VDD VSS N006 tl082
XU2 0 N011 VDD VSS N007 tl082
XU3 0 N013 VDD VSS N002 tl082
XU4 0 N015 VDD VSS N016 tl082
XU8 0 N012 VDD VSS N009 tl082

* MULTIPLIER
XU5 N001 0 ve N006 0 vdd N003 N003 0 vss MPY634
XU6 N001 0 ve N007 0 vdd N004 N004 0 vss MPY634
XU7 N002 0 ve N008 0 vdd N005 N005 0 vss MPY634

* SUPPLY
VDD vdd 0 {Vsup}
VSS 0 vss {Vsup}
VE ve 0 {Vsup}

V4 N014 0 {Vx4}
V1 N008 0 PULSE(-100m 100m 0 1n 1n 500u 1m)
+         AC 1 0

* ANALYSIS
.ac dec 101 50 10k
*.tran 60m
.step param Vx4 1 100 20

.end
